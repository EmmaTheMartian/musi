module interpreter

pub struct Trace {
pub:
	file   string
	source string
	line   int
	column int
}
