module musi
