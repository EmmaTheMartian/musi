module musi

pub type Value = string | int | f32
